
module simple_and 
        (
            //input
            a,
            b,
            // output
            c
        );

    //port definition
    input a;
    input b;

    output c;

    // design implementation
    
    assign c = a & b;

endmodule

    
